module();
endmodule
